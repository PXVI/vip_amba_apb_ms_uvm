// *******************************************************
// Date Created   : 31 May, 2019
// Author         : :P
// *******************************************************


