// ***********************************
// ************** :P *****************
// ***********************************
// Date Created : 21 May, 2019

`ifndef COMMON_TB_DEFINES_PARAMS
// Defines Section
// ---------------


// Parameter Section
// -----------------

`endif
