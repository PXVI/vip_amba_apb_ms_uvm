// *******************************************************
// Date Created   : 05 June, 2019
// Author         : :P
// *******************************************************

interface vip_amba_apb_bridge_bfm_interface `VIP_AMBA_APB_BRIDGE_DECL;

  // Interface Signals Declaration

endinterface
