// *******************************************************
// Date Created   : 01 June, 2019
// Author         : :P
// *******************************************************


