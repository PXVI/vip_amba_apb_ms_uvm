// *******************************************************
// Date Created   : 07 June, 2019
// Author         : :P
// *******************************************************

interface vip_amba_apb_slave_bfm_interface `VIP_AMBA_APB_SLAVE_DECL;

  // Interface Signal Declarations

endinterface
