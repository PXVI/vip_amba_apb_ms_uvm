// ***********************************
// ************** :P *****************
// ***********************************
// Date Created : 21 May, 2019

`ifndef COMMON_TB_DEFINES_PARAMS
// Defines Section
// ---------------

// Local Parameter Section
// -----------------------

`define VIP_AMBA_APB_SLAVE_PARAM				#( )

// -----------------------
`endif
